module ahb2apb();


endmodule
